// PLL.v

// Generated using ACDS version 13.0sp1 232 at 2019.04.16.02:32:59

`timescale 1 ps / 1 ps
module PLL (
		input  wire  clock_in_clk,  //  clock_in.clk
		input  wire  reset_reset,   //     reset.reset
		output wire  clock_out_clk  // clock_out.clk
	);

	PLL_altpll_0 altpll_0 (
		.clk       (clock_in_clk),  //       inclk_interface.clk
		.reset     (reset_reset),   // inclk_interface_reset.reset
		.read      (),              //             pll_slave.read
		.write     (),              //                      .write
		.address   (),              //                      .address
		.readdata  (),              //                      .readdata
		.writedata (),              //                      .writedata
		.c0        (clock_out_clk), //                    c0.clk
		.areset    (),              //        areset_conduit.export
		.locked    (),              //        locked_conduit.export
		.phasedone ()               //     phasedone_conduit.export
	);

endmodule
